module ACC (
	input Load, Sh, Ad, Clk, rst,
	input [8:0] Entradas,
	output [8:0] Saidas
);

	//Aqui entra a implementação do ckt

endmodule

