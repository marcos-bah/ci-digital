module counter (
    input clk, rst, ena,
    output reg ack,
    output reg [7:0] addr_bus
);
    
endmodule