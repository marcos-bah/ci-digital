module CONTROL (
	input Clk, K, St, M, rst,
	output Idle, Done, Load, Sh, Ad
);

	//Aqui entra a implementação do ckt

endmodule
