//! Módulo inversor da Aula 01
module inversor (
    input a, //! Entrada
    output b //! Saída
);
    assign b = ~a;
endmodule