module inversor (s, a);
output s;
input a;
  assign s = ~ a;
endmodule
