module Multiplicador_TB();




endmodule

