module Adder (
	input [3:0] OperandoA, OperandoB,
	output [4:0] Soma
);
//Aqui entra a implementação do ckt

endmodule

