module conversorA (
    input H,G,F,E,
    output A
);
    assign A = H;
endmodule