module portanou (s, a, b);

input a, b;
output s;

nor I1 (s, a, b);

endmodule
