module ieee754_adder_subtb;
    reg  [31:0] a;
    reg  [31:0] b;
    reg         op;
    wire [31:0] result;

    ieee754_adder_sub uut (
        .a(a),
        .b(b),
        .op(op),
        .result(result)
    );

    initial begin
        $monitor("Tempo=%0t | op=%b | a=%b | b=%b | result=%b", $time, op, a, b, result);

        a = 32'b0_10000001_00000000000000000000000; // 4.0
        b = 32'b0_01111111_00000000000000000000000; // 1.0
        op = 1; #10; // 4.0 + 1.0
        op = 0; #10; // 4.0 - 1.0

        a = 32'b1_10000000_00000000000000000000000; // -2.0
        b = 32'b0_01111111_00000000000000000000000; // 1.0
        op = 1; #10; // -2.0 + 1.0
        op = 0; #10; // -2.0 - 1.0

        a = 32'b0_10000000_00000000000000000000000; // 2.0
        b = 32'b0_10000000_00000000000000000000000; // 2.0
        op = 0; #10; // 2.0 - 2.0

        $stop;
    end

endmodule
