module ula (
    input ena, clk,
    input [3:0] op1, op2, op_sel,
    output reg [3:0] res,
    output reg ula_ack
);
    
endmodule