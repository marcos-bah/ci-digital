module Counter (
	input Load, Clk, rst,
	output K
);

	//Aqui entra a implementação do ckt

endmodule
