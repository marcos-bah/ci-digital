module topo (
    input clk, rst
);
    
endmodule