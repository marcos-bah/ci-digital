module somador_3bits_bcd_tb ();

reg [11:0] A, B;
reg C_in;
wire [11:0] out;
wire C_out;

somador_3bits_bcd somador (
    .A(A),
    .B(B),
    .Cin(C_in),
    .Cout(C_out),
    .Y(out)
);

initial begin
    $display("\n");
    $monitor("A: %b + B: %b + Cin: %b = Out: %b | C_out: %b", A, B, C_in, out, C_out);

    // 000 + 000 + 0 = 000
    A = 12'b0000_0000_0000;
    B = 12'b0000_0000_0000;
    C_in = 0;
    #10;

    // 001 + 002 + 0 = 003
    A = 12'b0000_0000_0001; // 001
    B = 12'b0000_0000_0010; // 002
    C_in = 0;
    #10;

    // 001 + 003 + 1 = 005
    A = 12'b0000_0000_0001; // 001
    B = 12'b0000_0000_0011; // 003
    C_in = 1;
    #10;

    // 010 + 004 + 0 = 014
    A = 12'b0000_0001_0000; // 010
    B = 12'b0000_0000_0100; // 004
    C_in = 0;
    #10;

    // 123 + 456 + 0 = 579
    A = 12'b0001_0010_0011; // 123
    B = 12'b0100_0101_0110; // 456
    C_in = 0;
    #10;

    // 999 + 001 + 0 = 1000 (overflow test)
    A = 12'b1001_1001_1001; // 999
    B = 12'b0000_0000_0001; // 001
    C_in = 0;
    #10;

    // 999 + 999 + 0 = 1998 (overflow test)
    A = 12'b1001_1001_1001; // 999
    B = 12'b1001_1001_1001; // 999
    C_in = 0;
    #10;
end
endmodule

