module mux16x1_tb();
    reg [15:0] in;
    reg [3:0] sel; 
    wire out;

    mux16x1 uut (.in(in), .sel(sel), .out(out));

    initial begin
        in = 16'b0101_0101_0101_0101;
        $display("\n");
        sel = 4'b0000; #10;
        sel = 4'b0001; #10;
        sel = 4'b0010; #10;
        sel = 4'b0011; #10;
        sel = 4'b0100; #10;
        sel = 4'b0101; #10;
        sel = 4'b0110; #10;
        sel = 4'b0111; #10;
    end

    initial begin
        $monitor("Tempo: %0t | Entrada: %b | Sel %b | Saída: %b", $time ,in, sel, out);
    end

endmodule